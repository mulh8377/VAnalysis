module tokenf

//to do
pub fn tokenize(expr string) [] string {
	res := []string
	return res
}